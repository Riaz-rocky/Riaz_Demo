riaz new git file
acvsjj