i want to understand check out command 