fhfhj
cvbd
ls
uu