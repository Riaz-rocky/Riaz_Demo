fhfhj
cvbd
riaz
ls
uu
