riaz new git file
acvsjj
jkd
