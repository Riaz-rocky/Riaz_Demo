riaz new git file