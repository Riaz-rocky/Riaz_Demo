fhfhj
cvbd
