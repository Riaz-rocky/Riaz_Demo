fhfhj
cvbd
riaz
riaz1
ls
uu
