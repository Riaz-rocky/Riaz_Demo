fhfhj
